library ieee;
use ieee.std_logic_1164.all;

-- This defines the data type state used in multiple files
package DataTypePackage is

	type state is (
						init,
						s0a,s0b,s0c,
						s1a,s1b,
						s2a,s2b,
						s3a,s3b,
						s4,
						s5a,s5b,
						s6a,s6b,
						s7a,s7b,s7c,
						s8a,s8b,
						s9a,s9b,s9c,
						s10a,s10b,
						s11,
						s12a,s12b,
						s13,
						s14a,s14b,
						s15,
						s16a,s16b,s16c,
						s17a,s17b,
						s18a,s18b,
						s19a,s19b
						);
						
end package;